library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Sbox is
    Port ( Byte_in : in STD_LOGIC_VECTOR (7 downto 0);
           Byte_out : out STD_LOGIC_VECTOR (7 downto 0));
end Sbox;

architecture Behavioral of Sbox is

begin
    Process(Byte_in)
        begin
            case Byte_in is
                when x"00" => Byte_out <= x"63";
                when x"01" => Byte_out <= x"7c";
                when x"02" => Byte_out <= x"77";
                when x"03" => Byte_out <= x"7b";
                when x"04" => Byte_out <= x"f2";
                when x"05" => Byte_out <= x"6b";
                when x"06" => Byte_out <= x"6f";
                when x"07" => Byte_out <= x"c5";
                when x"08" => Byte_out <= x"30";
                when x"09" => Byte_out <= x"01";
                when x"0a" => Byte_out <= x"67";
                when x"0b" => Byte_out <= x"2b";
                when x"0c" => Byte_out <= x"fe";
                when x"0d" => Byte_out <= x"d7";
                when x"0e" => Byte_out <= x"ab";
                when x"0f" => Byte_out <= x"76";
                when x"10" => Byte_out <= x"ca";
                when x"11" => Byte_out <= x"82";
                when x"12" => Byte_out <= x"c9";
                when x"13" => Byte_out <= x"7d";
                when x"14" => Byte_out <= x"fa";
                when x"15" => Byte_out <= x"59";
                when x"16" => Byte_out <= x"47";
                when x"17" => Byte_out <= x"f0";
                when x"18" => Byte_out <= x"ad";
                when x"19" => Byte_out <= x"d4";
                when x"1a" => Byte_out <= x"a2";
                when x"1b" => Byte_out <= x"af";
                when x"1c" => Byte_out <= x"9c";
                when x"1d" => Byte_out <= x"a4";
                when x"1e" => Byte_out <= x"72";
                when x"1f" => Byte_out <= x"c0";
                when x"20" => Byte_out <= x"b7";
                when x"21" => Byte_out <= x"fd";
                when x"22" => Byte_out <= x"93";
                when x"23" => Byte_out <= x"26";
                when x"24" => Byte_out <= x"36";
                when x"25" => Byte_out <= x"3f";
                when x"26" => Byte_out <= x"f7";
                when x"27" => Byte_out <= x"cc";
                when x"28" => Byte_out <= x"34";
                when x"29" => Byte_out <= x"a5";
                when x"2a" => Byte_out <= x"e5";
                when x"2b" => Byte_out <= x"f1";
                when x"2c" => Byte_out <= x"71";
                when x"2d" => Byte_out <= x"d8";
                when x"2e" => Byte_out <= x"31";
                when x"2f" => Byte_out <= x"15";
                when x"30" => Byte_out <= x"04";
                when x"31" => Byte_out <= x"c7";
                when x"32" => Byte_out <= x"23";
                when x"33" => Byte_out <= x"c3";
                when x"34" => Byte_out <= x"18";
                when x"35" => Byte_out <= x"96";
                when x"36" => Byte_out <= x"05";
                when x"37" => Byte_out <= x"9a";
                when x"38" => Byte_out <= x"07";
                when x"39" => Byte_out <= x"12";
                when x"3a" => Byte_out <= x"80";
                when x"3b" => Byte_out <= x"e2";
                when x"3c" => Byte_out <= x"eb";
                when x"3d" => Byte_out <= x"27";
                when x"3e" => Byte_out <= x"b2";
                when x"3f" => Byte_out <= x"75";
                when x"40" => Byte_out <= x"09";
                when x"41" => Byte_out <= x"83";
                when x"42" => Byte_out <= x"2c";
                when x"43" => Byte_out <= x"1a";
                when x"44" => Byte_out <= x"1b";
                when x"45" => Byte_out <= x"6e";
                when x"46" => Byte_out <= x"5a";
                when x"47" => Byte_out <= x"a0";
                when x"48" => Byte_out <= x"52";
                when x"49" => Byte_out <= x"3b";
                when x"4a" => Byte_out <= x"d6";
                when x"4b" => Byte_out <= x"b3";
                when x"4c" => Byte_out <= x"29";
                when x"4d" => Byte_out <= x"e3";
                when x"4e" => Byte_out <= x"2f";
                when x"4f" => Byte_out <= x"84";
                when x"50" => Byte_out <= x"53";
                when x"51" => Byte_out <= x"d1";
                when x"52" => Byte_out <= x"00";
                when x"53" => Byte_out <= x"ed";
                when x"54" => Byte_out <= x"20";
                when x"55" => Byte_out <= x"fc";
                when x"56" => Byte_out <= x"b1";
                when x"57" => Byte_out <= x"5b";
                when x"58" => Byte_out <= x"6a";
                when x"59" => Byte_out <= x"cb";
                when x"5a" => Byte_out <= x"be";
                when x"5b" => Byte_out <= x"39";
                when x"5c" => Byte_out <= x"4a";
                when x"5d" => Byte_out <= x"4c";
                when x"5e" => Byte_out <= x"58";
                when x"5f" => Byte_out <= x"cf";
                when x"60" => Byte_out <= x"d0";
                when x"61" => Byte_out <= x"ef";
                when x"62" => Byte_out <= x"aa";
                when x"63" => Byte_out <= x"fb";
                when x"64" => Byte_out <= x"43";
                when x"65" => Byte_out <= x"4d";
                when x"66" => Byte_out <= x"33";
                when x"67" => Byte_out <= x"85";
                when x"68" => Byte_out <= x"45";
                when x"69" => Byte_out <= x"f9";
                when x"6a" => Byte_out <= x"02";
                when x"6b" => Byte_out <= x"7f";
                when x"6c" => Byte_out <= x"50";
                when x"6d" => Byte_out <= x"3c";
                when x"6e" => Byte_out <= x"9f";
                when x"6f" => Byte_out <= x"a8";
                when x"70" => Byte_out <= x"51";
                when x"71" => Byte_out <= x"a3";
                when x"72" => Byte_out <= x"40";
                when x"73" => Byte_out <= x"8f";
                when x"74" => Byte_out <= x"92";
                when x"75" => Byte_out <= x"9d";
                when x"76" => Byte_out <= x"38";
                when x"77" => Byte_out <= x"f5";
                when x"78" => Byte_out <= x"bc";
                when x"79" => Byte_out <= x"b6";
                when x"7a" => Byte_out <= x"da";
                when x"7b" => Byte_out <= x"21";
                when x"7c" => Byte_out <= x"10";
                when x"7d" => Byte_out <= x"ff";
                when x"7e" => Byte_out <= x"f3";
                when x"7f" => Byte_out <= x"d2";
                when x"80" => Byte_out <= x"cd";
                when x"81" => Byte_out <= x"0c";
                when x"82" => Byte_out <= x"13";
                when x"83" => Byte_out <= x"ec";
                when x"84" => Byte_out <= x"5f";
                when x"85" => Byte_out <= x"97";
                when x"86" => Byte_out <= x"44";
                when x"87" => Byte_out <= x"17";
                when x"88" => Byte_out <= x"c4";
                when x"89" => Byte_out <= x"a7";
                when x"8a" => Byte_out <= x"7e";
                when x"8b" => Byte_out <= x"3d";
                when x"8c" => Byte_out <= x"64";
                when x"8d" => Byte_out <= x"5d";
                when x"8e" => Byte_out <= x"19";
                when x"8f" => Byte_out <= x"73";
                when x"90" => Byte_out <= x"60";
                when x"91" => Byte_out <= x"81";
                when x"92" => Byte_out <= x"4f";
                when x"93" => Byte_out <= x"dc";
                when x"94" => Byte_out <= x"22";
                when x"95" => Byte_out <= x"2a";
                when x"96" => Byte_out <= x"90";
                when x"97" => Byte_out <= x"88";
                when x"98" => Byte_out <= x"46";
                when x"99" => Byte_out <= x"ee";
                when x"9a" => Byte_out <= x"b8";
                when x"9b" => Byte_out <= x"14";
                when x"9c" => Byte_out <= x"de";
                when x"9d" => Byte_out <= x"5e";
                when x"9e" => Byte_out <= x"0b";
                when x"9f" => Byte_out <= x"db";
                when x"a0" => Byte_out <= x"e0";
                when x"a1" => Byte_out <= x"32";
                when x"a2" => Byte_out <= x"3a";
                when x"a3" => Byte_out <= x"0a";
                when x"a4" => Byte_out <= x"49";
                when x"a5" => Byte_out <= x"06";
                when x"a6" => Byte_out <= x"24";
                when x"a7" => Byte_out <= x"5c";
                when x"a8" => Byte_out <= x"c2";
                when x"a9" => Byte_out <= x"d3";
                when x"aa" => Byte_out <= x"ac";
                when x"ab" => Byte_out <= x"62";
                when x"ac" => Byte_out <= x"91";
                when x"ad" => Byte_out <= x"95";
                when x"ae" => Byte_out <= x"e4";
                when x"af" => Byte_out <= x"79";
                when x"b0" => Byte_out <= x"e7";
                when x"b1" => Byte_out <= x"c8";
                when x"b2" => Byte_out <= x"37";
                when x"b3" => Byte_out <= x"6d";
                when x"b4" => Byte_out <= x"8d";
                when x"b5" => Byte_out <= x"d5";
                when x"b6" => Byte_out <= x"4e";
                when x"b7" => Byte_out <= x"a9";
                when x"b8" => Byte_out <= x"6c";
                when x"b9" => Byte_out <= x"56";
                when x"ba" => Byte_out <= x"f4";
                when x"bb" => Byte_out <= x"ea";
                when x"bc" => Byte_out <= x"65";
                when x"bd" => Byte_out <= x"7a";
                when x"be" => Byte_out <= x"ae";
                when x"bf" => Byte_out <= x"08";
                when x"c0" => Byte_out <= x"ba";
                when x"c1" => Byte_out <= x"78";
                when x"c2" => Byte_out <= x"25";
                when x"c3" => Byte_out <= x"2e";
                when x"c4" => Byte_out <= x"1c";
                when x"c5" => Byte_out <= x"a6";
                when x"c6" => Byte_out <= x"b4";
                when x"c7" => Byte_out <= x"c6";
                when x"c8" => Byte_out <= x"e8";
                when x"c9" => Byte_out <= x"dd";
                when x"ca" => Byte_out <= x"74";
                when x"cb" => Byte_out <= x"1f";
                when x"cc" => Byte_out <= x"4b";
                when x"cd" => Byte_out <= x"bd";
                when x"ce" => Byte_out <= x"8b";
                when x"cf" => Byte_out <= x"8a";
                when x"d0" => Byte_out <= x"70";
                when x"d1" => Byte_out <= x"3e";
                when x"d2" => Byte_out <= x"b5";
                when x"d3" => Byte_out <= x"66";
                when x"d4" => Byte_out <= x"48";
                when x"d5" => Byte_out <= x"03";
                when x"d6" => Byte_out <= x"f6";
                when x"d7" => Byte_out <= x"0e";
                when x"d8" => Byte_out <= x"61";
                when x"d9" => Byte_out <= x"35";
                when x"da" => Byte_out <= x"57";
                when x"db" => Byte_out <= x"b9";
                when x"dc" => Byte_out <= x"86";
                when x"dd" => Byte_out <= x"c1";
                when x"de" => Byte_out <= x"1d";
                when x"df" => Byte_out <= x"9e";
                when x"e0" => Byte_out <= x"e1";
                when x"e1" => Byte_out <= x"f8";
                when x"e2" => Byte_out <= x"98";
                when x"e3" => Byte_out <= x"11";
                when x"e4" => Byte_out <= x"69";
                when x"e5" => Byte_out <= x"d9";
                when x"e6" => Byte_out <= x"8e";
                when x"e7" => Byte_out <= x"94";
                when x"e8" => Byte_out <= x"9b";
                when x"e9" => Byte_out <= x"1e";
                when x"ea" => Byte_out <= x"87";
                when x"eb" => Byte_out <= x"e9";
                when x"ec" => Byte_out <= x"ce";
                when x"ed" => Byte_out <= x"55";
                when x"ee" => Byte_out <= x"28";
                when x"ef" => Byte_out <= x"df";
                when x"f0" => Byte_out <= x"8c";
                when x"f1" => Byte_out <= x"a1";
                when x"f2" => Byte_out <= x"89";
                when x"f3" => Byte_out <= x"0d";
                when x"f4" => Byte_out <= x"bf";
                when x"f5" => Byte_out <= x"e6";
                when x"f6" => Byte_out <= x"42";
                when x"f7" => Byte_out <= x"68";
                when x"f8" => Byte_out <= x"41";
                when x"f9" => Byte_out <= x"99";
                when x"fa" => Byte_out <= x"2d";
                when x"fb" => Byte_out <= x"0f";
                when x"fc" => Byte_out <= x"b0";
                when x"fd" => Byte_out <= x"54";
                when x"fe" => Byte_out <= x"bb";
                when x"ff" => Byte_out <= x"16";
                when others => Byte_out <= x"00";               
            end case;
    end Process;
    
end Behavioral;
